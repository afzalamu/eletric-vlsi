*** SPICE deck for cell inv_sim{lay} from library inv_20_10
*** Created on Thu Aug 17, 2023 12:04:27
*** Last revised on Thu Aug 17, 2023 12:20:17
*** Written on Thu Aug 17, 2023 17:39:18 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT inv_20_10__inv_20_10 FROM CELL inv_20_10{lay}
.SUBCKT inv_20_10__inv_20_10 gnd IN OUT vdd
Mnmos@0 OUT IN gnd gnd NMOS L=0.6U W=3U AS=16.2P AD=10.8P PS=25.8U PD=13.8U
Mpmos@0 OUT IN vdd vdd PMOS L=0.6U W=6U AS=23.4P AD=10.8P PS=31.8U PD=13.8U
.ENDS inv_20_10__inv_20_10

*** TOP LEVEL CELL: inv_sim{lay}
Xinv_20_1@0 gnd IN OUT vdd inv_20_10__inv_20_10

* Spice Code nodes in cell cell 'inv_sim{lay}'
vdd vdd 0 DC 5
vin in 0 DC 0
.dc vin 0 5 1m
.include "C:\ELECTRIC VLSI\C50.txt"
.END
